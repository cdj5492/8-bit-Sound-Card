-- Copyright (C) 2021  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.0 Build 842 10/21/2021 SJ Lite Edition"
-- CREATED		"Sat Mar  5 16:28:34 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Envelope IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		Ev1 :  IN  STD_LOGIC;
		Ev2 :  IN  STD_LOGIC;
		Ev3 :  IN  STD_LOGIC;
		Ev4 :  IN  STD_LOGIC;
		EvStore :  IN  STD_LOGIC;
		SetStartFlag :  IN  STD_LOGIC;
		LoopFlag :  IN  STD_LOGIC;
		ConstantVolumeFlag :  IN  STD_LOGIC;
		Env_Out :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END Envelope;

ARCHITECTURE bdf_type OF Envelope IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \4count_0\
	PORT(LDN : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 SETN : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \4count_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \4count_0\: COMPONENT IS true;

COMPONENT \4count_1\
	PORT(LDN : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 SETN : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC;
		 QD : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \4count_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \4count_1\: COMPONENT IS true;

COMPONENT busmux_2
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_2: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_2: COMPONENT IS true;

SIGNAL	Decay :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	Delay :  STD_LOGIC_VECTOR(3 TO 3);
SIGNAL	Env :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	DFF_inst18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	DFF_inst8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_44 <= '1';
SYNTHESIZED_WIRE_49 <= '1';
SYNTHESIZED_WIRE_51 <= '0';
SYNTHESIZED_WIRE_52 <= '1';
SYNTHESIZED_WIRE_18 <= '0';
SYNTHESIZED_WIRE_19 <= '1';
SYNTHESIZED_WIRE_54 <= '0';
SYNTHESIZED_WIRE_55 <= '1';
SYNTHESIZED_WIRE_34 <= '0';
SYNTHESIZED_WIRE_36 <= '1';
SYNTHESIZED_WIRE_38 <= '1';
SYNTHESIZED_WIRE_39 <= '1';
SYNTHESIZED_WIRE_40 <= '0';
SYNTHESIZED_WIRE_41 <= '1';




b2v_DecayC : 4count_0
PORT MAP(LDN => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_44,
		 A => SYNTHESIZED_WIRE_44,
		 D => SYNTHESIZED_WIRE_44,
		 CIN => SYNTHESIZED_WIRE_44,
		 DNUP => SYNTHESIZED_WIRE_44,
		 CLK => SYNTHESIZED_WIRE_45,
		 SETN => SYNTHESIZED_WIRE_44,
		 C => SYNTHESIZED_WIRE_44,
		 CLRN => SYNTHESIZED_WIRE_44,
		 QA => Decay(0),
		 QB => Decay(1),
		 QC => Decay(2));


b2v_Divider : 4count_1
PORT MAP(LDN => SYNTHESIZED_WIRE_9,
		 B => SYNTHESIZED_WIRE_46,
		 A => SYNTHESIZED_WIRE_47,
		 D => SYNTHESIZED_WIRE_48,
		 CIN => SYNTHESIZED_WIRE_49,
		 DNUP => SYNTHESIZED_WIRE_49,
		 CLK => CLK,
		 SETN => SYNTHESIZED_WIRE_49,
		 C => SYNTHESIZED_WIRE_50,
		 CLRN => SYNTHESIZED_WIRE_49,
		 QA => SYNTHESIZED_WIRE_26,
		 QB => SYNTHESIZED_WIRE_28,
		 QC => SYNTHESIZED_WIRE_27,
		 QD => SYNTHESIZED_WIRE_29);


b2v_inst : busmux_2
PORT MAP(sel => DFF_inst18,
		 dataa => Decay,
		 datab => Env,
		 result => Env_Out);


PROCESS(EvStore,SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_50 <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	SYNTHESIZED_WIRE_50 <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	SYNTHESIZED_WIRE_50 <= Ev3;
END IF;
END PROCESS;





SYNTHESIZED_WIRE_37 <= NOT(CLK AND SYNTHESIZED_WIRE_53);


SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_53 AND DFF_inst8);


PROCESS(EvStore,SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_47 <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	SYNTHESIZED_WIRE_47 <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	SYNTHESIZED_WIRE_47 <= Ev1;
END IF;
END PROCESS;




PROCESS(CLK,SYNTHESIZED_WIRE_18,SYNTHESIZED_WIRE_19)
BEGIN
IF (SYNTHESIZED_WIRE_18 = '0') THEN
	DFF_inst18 <= '0';
ELSIF (SYNTHESIZED_WIRE_19 = '0') THEN
	DFF_inst18 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst18 <= ConstantVolumeFlag;
END IF;
END PROCESS;



PROCESS(EvStore,SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	SYNTHESIZED_WIRE_46 <= Ev2;
END IF;
END PROCESS;







PROCESS(EvStore,SYNTHESIZED_WIRE_54,SYNTHESIZED_WIRE_55)
BEGIN
IF (SYNTHESIZED_WIRE_54 = '0') THEN
	Env(0) <= '0';
ELSIF (SYNTHESIZED_WIRE_55 = '0') THEN
	Env(0) <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	Env(0) <= SYNTHESIZED_WIRE_47;
END IF;
END PROCESS;


PROCESS(EvStore,SYNTHESIZED_WIRE_54,SYNTHESIZED_WIRE_55)
BEGIN
IF (SYNTHESIZED_WIRE_54 = '0') THEN
	Env(3) <= '0';
ELSIF (SYNTHESIZED_WIRE_55 = '0') THEN
	Env(3) <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	Env(3) <= SYNTHESIZED_WIRE_48;
END IF;
END PROCESS;




SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_45);



SYNTHESIZED_WIRE_35 <= NOT(SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27 OR SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29);


PROCESS(EvStore,SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_48 <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	SYNTHESIZED_WIRE_48 <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	SYNTHESIZED_WIRE_48 <= Ev4;
END IF;
END PROCESS;


PROCESS(EvStore,SYNTHESIZED_WIRE_54,SYNTHESIZED_WIRE_55)
BEGIN
IF (SYNTHESIZED_WIRE_54 = '0') THEN
	Env(2) <= '0';
ELSIF (SYNTHESIZED_WIRE_55 = '0') THEN
	Env(2) <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	Env(2) <= SYNTHESIZED_WIRE_50;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_36)
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	SYNTHESIZED_WIRE_45 <= '0';
ELSIF (SYNTHESIZED_WIRE_36 = '0') THEN
	SYNTHESIZED_WIRE_45 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_45 <= SYNTHESIZED_WIRE_35;
END IF;
END PROCESS;


PROCESS(SetStartFlag,SYNTHESIZED_WIRE_37,SYNTHESIZED_WIRE_39)
BEGIN
IF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_53 <= '0';
ELSIF (SYNTHESIZED_WIRE_39 = '0') THEN
	SYNTHESIZED_WIRE_53 <= '1';
ELSIF (RISING_EDGE(SetStartFlag)) THEN
	SYNTHESIZED_WIRE_53 <= SYNTHESIZED_WIRE_38;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_40,SYNTHESIZED_WIRE_41)
BEGIN
IF (SYNTHESIZED_WIRE_40 = '0') THEN
	DFF_inst8 <= '0';
ELSIF (SYNTHESIZED_WIRE_41 = '0') THEN
	DFF_inst8 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst8 <= LoopFlag;
END IF;
END PROCESS;


PROCESS(EvStore,SYNTHESIZED_WIRE_54,SYNTHESIZED_WIRE_55)
BEGIN
IF (SYNTHESIZED_WIRE_54 = '0') THEN
	Env(1) <= '0';
ELSIF (SYNTHESIZED_WIRE_55 = '0') THEN
	Env(1) <= '1';
ELSIF (RISING_EDGE(EvStore)) THEN
	Env(1) <= SYNTHESIZED_WIRE_46;
END IF;
END PROCESS;


END bdf_type;