-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sat Mar 05 19:03:33 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Envelope IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		EvStore :  IN  STD_LOGIC;
		SetStartFlag :  IN  STD_LOGIC;
		LoopFlag :  IN  STD_LOGIC;
		ConstantVolumeFlag :  IN  STD_LOGIC;
		Ev3t :  IN  STD_LOGIC;
		Ev2t :  IN  STD_LOGIC;
		Ev1t :  IN  STD_LOGIC;
		Ev4t :  IN  STD_LOGIC;
		tstIn :  IN  STD_LOGIC;
		tstOut :  OUT  STD_LOGIC;
		Env_Out :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END Envelope;

ARCHITECTURE bdf_type OF Envelope IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \4count_0\
	PORT(LDN : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 SETN : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \4count_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \4count_0\: COMPONENT IS true;

COMPONENT \4count_1\
	PORT(LDN : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 SETN : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC;
		 QD : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \4count_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \4count_1\: COMPONENT IS true;

COMPONENT busmux_2
	PORT(sel : IN STD_LOGIC;
		 dataa : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 datab : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COMPONENT;
ATTRIBUTE black_box OF busmux_2: COMPONENT IS true;
ATTRIBUTE noopt OF busmux_2: COMPONENT IS true;

SIGNAL	Decay :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	Delay :  STD_LOGIC_VECTOR(3 TO 3);
SIGNAL	EV :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	DFF_inst8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	DFF_inst18 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_45 <= '1';
SYNTHESIZED_WIRE_47 <= '1';
SYNTHESIZED_WIRE_50 <= '0';
SYNTHESIZED_WIRE_52 <= '1';
SYNTHESIZED_WIRE_22 <= '1';
SYNTHESIZED_WIRE_24 <= '1';
SYNTHESIZED_WIRE_35 <= '1';
SYNTHESIZED_WIRE_38 <= '1';
SYNTHESIZED_WIRE_40 <= '1';
SYNTHESIZED_WIRE_41 <= '1';
SYNTHESIZED_WIRE_42 <= '0';
SYNTHESIZED_WIRE_44 <= '1';




b2v_DecayC : 4count_0
PORT MAP(LDN => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_45,
		 A => SYNTHESIZED_WIRE_45,
		 D => SYNTHESIZED_WIRE_45,
		 CIN => SYNTHESIZED_WIRE_45,
		 DNUP => SYNTHESIZED_WIRE_45,
		 CLK => SYNTHESIZED_WIRE_46,
		 SETN => SYNTHESIZED_WIRE_45,
		 C => SYNTHESIZED_WIRE_45,
		 CLRN => SYNTHESIZED_WIRE_45,
		 QA => Decay(0),
		 QB => Decay(1),
		 QC => Decay(2));


b2v_Divider : 4count_1
PORT MAP(LDN => SYNTHESIZED_WIRE_9,
		 B => EV(1),
		 A => EV(0),
		 D => EV(3),
		 CIN => SYNTHESIZED_WIRE_47,
		 DNUP => SYNTHESIZED_WIRE_47,
		 CLK => SYNTHESIZED_WIRE_48,
		 SETN => SYNTHESIZED_WIRE_47,
		 C => EV(2),
		 CLRN => SYNTHESIZED_WIRE_47,
		 QA => SYNTHESIZED_WIRE_28,
		 QB => SYNTHESIZED_WIRE_30,
		 QC => SYNTHESIZED_WIRE_29,
		 QD => SYNTHESIZED_WIRE_31);


SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_46 OR SYNTHESIZED_WIRE_49);


PROCESS(SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_50,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_50 = '0') THEN
	EV(2) <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	EV(2) <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_51)) THEN
	EV(2) <= Ev3t;
END IF;
END PROCESS;



tstOut <= NOT(tstIn);





SYNTHESIZED_WIRE_39 <= NOT(SYNTHESIZED_WIRE_48 AND SYNTHESIZED_WIRE_49);


SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_49 AND DFF_inst8);


PROCESS(SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_50,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_50 = '0') THEN
	EV(0) <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	EV(0) <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_51)) THEN
	EV(0) <= Ev1t;
END IF;
END PROCESS;




PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_22,SYNTHESIZED_WIRE_24)
BEGIN
IF (SYNTHESIZED_WIRE_22 = '0') THEN
	DFF_inst18 <= '0';
ELSIF (SYNTHESIZED_WIRE_24 = '0') THEN
	DFF_inst18 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_48)) THEN
	DFF_inst18 <= ConstantVolumeFlag;
END IF;
END PROCESS;



PROCESS(SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_50,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_50 = '0') THEN
	EV(1) <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	EV(1) <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_51)) THEN
	EV(1) <= Ev2t;
END IF;
END PROCESS;







SYNTHESIZED_WIRE_37 <= NOT(SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29 OR SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_31);


PROCESS(SYNTHESIZED_WIRE_51,SYNTHESIZED_WIRE_50,SYNTHESIZED_WIRE_52)
BEGIN
IF (SYNTHESIZED_WIRE_50 = '0') THEN
	EV(3) <= '0';
ELSIF (SYNTHESIZED_WIRE_52 = '0') THEN
	EV(3) <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_51)) THEN
	EV(3) <= Ev4t;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_51 <= NOT(EvStore);



PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_35,SYNTHESIZED_WIRE_38)
BEGIN
IF (SYNTHESIZED_WIRE_35 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_48)) THEN
	SYNTHESIZED_WIRE_46 <= SYNTHESIZED_WIRE_37;
END IF;
END PROCESS;


PROCESS(SetStartFlag,SYNTHESIZED_WIRE_39,SYNTHESIZED_WIRE_41)
BEGIN
IF (SYNTHESIZED_WIRE_39 = '0') THEN
	SYNTHESIZED_WIRE_49 <= '0';
ELSIF (SYNTHESIZED_WIRE_41 = '0') THEN
	SYNTHESIZED_WIRE_49 <= '1';
ELSIF (RISING_EDGE(SetStartFlag)) THEN
	SYNTHESIZED_WIRE_49 <= SYNTHESIZED_WIRE_40;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_48,SYNTHESIZED_WIRE_42,SYNTHESIZED_WIRE_44)
BEGIN
IF (SYNTHESIZED_WIRE_42 = '0') THEN
	DFF_inst8 <= '0';
ELSIF (SYNTHESIZED_WIRE_44 = '0') THEN
	DFF_inst8 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_48)) THEN
	DFF_inst8 <= LoopFlag;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_48 <= NOT(CLK);



b2v_insts : busmux_2
PORT MAP(sel => DFF_inst18,
		 dataa => Decay,
		 datab => EV,
		 result => Env_Out);


END bdf_type;